`timescale 1ns / 1ps

module tb_conv_top;

    localparam WT_DEPTH        = 4096;
    localparam WT_ADDR_WIDTH   = $clog2(WT_DEPTH);
    localparam BIAS_DEPTH      = 256;
    localparam BIAS_GROUP_BITS = $clog2(BIAS_DEPTH) - 1;
    localparam WT_LATENCY      = 3;
    localparam CONV_PE_PIPE    = 3;
    localparam PIPE_DEPTH      = WT_LATENCY + CONV_PE_PIPE + 1; // 7

    // ── DUT signals ──
    logic        clk, rst;

    logic [9:0]                    cfg_ci_groups;
    logic [BIAS_GROUP_BITS-1:0]    cfg_output_group;
    logic [WT_ADDR_WIDTH-1:0]      cfg_wt_base_addr;
    logic [15:0]                   cfg_in_channels;
    logic [15:0]                   cfg_img_width;
    logic                          cfg_use_maxpool;
    logic                          cfg_stride_2;
    logic [31:0]                   cfg_quant_m;
    logic [4:0]                    cfg_quant_n;
    logic                          cfg_use_relu;
    logic                          go;
    logic                          busy, done;

    logic                          bias_wr_en;
    logic [127:0]                  bias_wr_data;
    logic                          bias_wr_addr_rst;

    logic                          wt_wr_en;
    logic [71:0]                   wt_wr_data;
    logic                          wt_wr_addr_rst;

    logic [63:0]                   pixel_in;
    logic                          pixel_in_valid;
    logic                          pixel_in_last;

    logic [63:0]                   data_out;
    logic                          data_out_valid;

    // Debug
    logic [31:0]                   dbg_bias_out [0:7];
    logic                          dbg_bias_valid;
    logic [575:0]                  dbg_wt_data_out [0:7];
    logic                          dbg_wt_data_ready;
    logic                          dbg_conv_valid_in;
    logic                          dbg_conv_last_channel;
    logic [63:0]                   dbg_pixel_d2 [0:2][0:2];

    // ── DUT ──
    conv_top #(
        .WT_DEPTH   (WT_DEPTH),
        .BIAS_DEPTH (BIAS_DEPTH),
        .WT_LATENCY (WT_LATENCY),
        .CONV_PE_PIPE(CONV_PE_PIPE)
    ) u_dut (
        .clk(clk),
        .rst(rst),
        .cfg_ci_groups(cfg_ci_groups),
        .cfg_output_group(cfg_output_group),
        .cfg_wt_base_addr(cfg_wt_base_addr),
        .cfg_in_channels(cfg_in_channels),
        .cfg_img_width(cfg_img_width),
        .cfg_use_maxpool(cfg_use_maxpool),
        .cfg_stride_2(cfg_stride_2),
        .cfg_quant_m(cfg_quant_m),
        .cfg_quant_n(cfg_quant_n),
        .cfg_use_relu(cfg_use_relu),
        .go(go),
        .busy(busy),
        .done(done),
        .bias_wr_en(bias_wr_en),
        .bias_wr_data(bias_wr_data),
        .bias_wr_addr_rst(bias_wr_addr_rst),
        .wt_wr_en(wt_wr_en),
        .wt_wr_data(wt_wr_data),
        .wt_wr_addr_rst(wt_wr_addr_rst),
        .pixel_in(pixel_in),
        .pixel_in_valid(pixel_in_valid),
        .pixel_in_last(pixel_in_last),
        .data_out(data_out),
        .data_out_valid(data_out_valid),
        .dbg_bias_out(dbg_bias_out),
        .dbg_bias_valid(dbg_bias_valid),
        .dbg_wt_data_out(dbg_wt_data_out),
        .dbg_wt_data_ready(dbg_wt_data_ready),
        .dbg_conv_valid_in(dbg_conv_valid_in),
        .dbg_conv_last_channel(dbg_conv_last_channel),
        .dbg_pixel_d2(dbg_pixel_d2)
    );

    // ── Clock ──
    initial clk = 0;
    always #5 clk = ~clk; // 100 MHz

    // ── Timeout ──
    initial begin
        #5ms;
        $display("[%0t] TIMEOUT", $time);
        $finish;
    end

    int errors = 0;

    // ── pixel_at_pe: 1-cycle capture of dbg_pixel_d2 ──
    logic [63:0] pixel_at_pe [0:2][0:2];
    always_ff @(posedge clk) begin
        for (int r = 0; r < 3; r++)
            for (int c = 0; c < 3; c++)
                pixel_at_pe[r][c] <= dbg_pixel_d2[r][c];
    end

    // ═══════════════════════════════════════════════════════════
    //  Helpers
    // ═══════════════════════════════════════════════════════════

    task automatic reset_all();
        rst              = 1;
        go               = 0;
        cfg_ci_groups    = 0;
        cfg_output_group = 0;
        cfg_wt_base_addr = 0;
        cfg_in_channels  = 0;
        cfg_img_width    = 0;
        cfg_use_maxpool  = 0;
        cfg_stride_2     = 0;
        cfg_quant_m      = 0;
        cfg_quant_n      = 0;
        cfg_use_relu     = 0;
        bias_wr_en       = 0;
        bias_wr_data     = 0;
        bias_wr_addr_rst = 0;
        wt_wr_en         = 0;
        wt_wr_data       = 0;
        wt_wr_addr_rst   = 0;
        pixel_in         = 0;
        pixel_in_valid   = 0;
        pixel_in_last    = 0;
        repeat(5) @(posedge clk);
        rst = 0;
        repeat(2) @(posedge clk);
    endtask

    // Stream image pixels to Input DMA interface
    task automatic stream_image(input int img_w, input int img_h, input int ci_groups);
        for (int r = 0; r < img_h; r++) begin
            for (int c = 0; c < img_w; c++) begin
                for (int ci = 0; ci < ci_groups; ci++) begin
                    @(posedge clk);
                    pixel_in_valid <= 1;
                    // Pattern: {8 bits row, 8 bits col, 8 bits ci_group, repeated}
                    pixel_in       <= {2{8'(r), 8'(c), 8'(ci), 8'hAA}};
                    pixel_in_last  <= (r == img_h-1 && c == img_w-1 && ci == ci_groups-1);
                end
            end
        end
        @(posedge clk);
        pixel_in_valid <= 0;
        pixel_in_last  <= 0;
    endtask

    // Load 8 biases
    task automatic load_biases(input logic [31:0] b [0:7]);
        @(posedge clk);
        bias_wr_addr_rst <= 1;
        @(posedge clk);
        bias_wr_addr_rst <= 0;
        @(posedge clk);
        bias_wr_en   <= 1;
        bias_wr_data <= {b[3], b[2], b[1], b[0]};
        @(posedge clk);
        bias_wr_data <= {b[7], b[6], b[5], b[4]};
        @(posedge clk);
        bias_wr_en   <= 0;
    endtask

    // Load weights
    task automatic load_weights(input int ci_groups, input logic [7:0] wt_val);
        logic [71:0] wt_word = {9{wt_val}};
        @(posedge clk);
        wt_wr_addr_rst <= 1;
        @(posedge clk);
        wt_wr_addr_rst <= 0;
        for (int addr = 0; addr < ci_groups; addr++) begin
            for (int bank = 0; bank < 8; bank++) begin
                for (int uram = 0; uram < 8; uram++) begin
                    @(posedge clk);
                    wt_wr_en   <= 1;
                    wt_wr_data <= wt_word;
                end
            end
        end
        @(posedge clk);
        wt_wr_en <= 0;
    endtask

    task automatic pulse_go();
        @(posedge clk);
        go <= 1;
        @(posedge clk);
        go <= 0;
    endtask

    task automatic wait_done(input int max_cycles);
        for (int i = 0; i < max_cycles; i++) begin
            @(posedge clk);
            if (done) return;
        end
        $display("[%0t] ERROR: done not asserted within %0d cycles", $time, max_cycles);
        errors++;
    endtask

    // ═══════════════════════════════════════════════════════════
    //  Tests
    // ═══════════════════════════════════════════════════════════

    task automatic test_kernel_window();
        $display("\n=== Test 1: Kernel Window + Pixel Delay ===");
        cfg_img_width   = 16'd4;
        cfg_in_channels = 16'd8;
        cfg_ci_groups   = 10'd1;
        fork
            stream_image(4, 4, 1);
            begin
                int timeout = 0;
                while (dbg_pixel_d2[1][1] == 0 && timeout < 100) begin
                    @(posedge clk);
                    timeout++;
                end
                if (timeout >= 100) begin
                    $display("  ERROR: No data reached pixel_d2");
                    errors++;
                end else begin
                    $display("  Data reached pixel_d2 at cycle %0d", timeout);
                end
            end
        join
        $display("  Test 1 done");
    endtask

    task automatic test_bias_load();
        logic [31:0] test_biases [0:7];
        $display("\n=== Test 2: Bias loading + readback ===");
        test_biases = '{32'd10, 32'd20, 32'd30, 32'd40, 32'd50, 32'd60, 32'd70, 32'd80};
        load_biases(test_biases);
        cfg_ci_groups    = 10'd1;
        cfg_output_group = 7'd0;
        cfg_wt_base_addr = 12'd0;
        cfg_img_width    = 16'd4;
        cfg_in_channels  = 16'd8;
        pulse_go();
        wait(dbg_bias_valid);
        @(negedge clk);
        for (int i = 0; i < 8; i++) begin
            if (dbg_bias_out[i] !== test_biases[i]) begin
                $display("  ERROR: bias_out[%0d] = %0d, expected %0d", i, dbg_bias_out[i], test_biases[i]);
                errors++;
            end
        end
        stream_image(4, 4, 1);
        wait_done(100);
        $display("  Test 2 done");
    endtask

    task automatic test_pipeline_timing();
        localparam CI_GROUPS = 1;
        int valid_count = 0;
        $display("\n=== Test 3: Pipeline timing (ci_groups=1, 4x4 image) ===");
        load_biases('{default: 32'd0});
        load_weights(CI_GROUPS, 8'd1);
        cfg_ci_groups    = CI_GROUPS;
        cfg_output_group = 7'd0;
        cfg_wt_base_addr = 12'd0;
        cfg_img_width    = 16'd4;
        cfg_in_channels  = 16'd8;
        pulse_go();
        fork
            stream_image(4, 4, CI_GROUPS);
            begin
                while (!done) begin
                    @(negedge clk);
                    if (dbg_conv_valid_in) begin
                        valid_count++;
                        if (!dbg_wt_data_ready) begin
                            $display("  ERROR: conv_valid_in but !wt_data_ready");
                            errors++;
                        end
                    end
                end
            end
        join
        // 4x4 image, 3x3 kernel -> 2x2 windows
        if (valid_count !== 4) begin
            $display("  ERROR: expected 4 conv_valid_in, got %0d", valid_count);
            errors++;
        end
        $display("  Test 3 done");
    endtask

    task automatic test_multi_ci();
        localparam CI_GROUPS = 2;
        int valid_count = 0;
        int last_ch_count = 0;
        $display("\n=== Test 4: Multi ci_groups=2, 4x4 image ===");
        load_biases('{default: 32'd0});
        load_weights(CI_GROUPS, 8'd1);
        cfg_ci_groups    = CI_GROUPS;
        cfg_output_group = 7'd0;
        cfg_wt_base_addr = 12'd0;
        cfg_img_width    = 16'd4;
        cfg_in_channels  = 16'd16;
        pulse_go();
        fork
            stream_image(4, 4, CI_GROUPS);
            begin
                while (!done) begin
                    @(negedge clk);
                    if (dbg_conv_valid_in) begin
                        valid_count++;
                        if (dbg_conv_last_channel) last_ch_count++;
                    end
                end
            end
        join
        if (valid_count !== 8) begin
            $display("  ERROR: expected 8 conv_valid_in, got %0d", valid_count);
            errors++;
        end
        if (last_ch_count !== 4) begin
            $display("  ERROR: expected 4 last_channel, got %0d", last_ch_count);
            errors++;
        end
        $display("  Test 4 done");
    endtask

    initial begin
        $dumpfile("tb_conv_top.vcd");
        $dumpvars(0, tb_conv_top);
        reset_all();
        test_kernel_window();
        reset_all();
        test_bias_load();
        reset_all();
        test_pipeline_timing();
        reset_all();
        test_multi_ci();
        #100;
        $display("\n════════════════════════════════════");
        if (errors == 0) $display("ALL TESTS PASSED");
        else $display("FAILED with %0d errors", errors);
        $display("════════════════════════════════════\n");
        $finish;
    end

endmodule
