module delayLine #(
    parameter WIDTH = 64,
    parameter MAX_DEPTH = 128
)(
    input logic clk,
    input logic rst,
    input logic en,
    input logic [7:0] delay_depth,// Cin/8
    input logic [WIDTH-1:0] din,
    output logic [WIDTH-1:0] dout
);

(* ram_style = "distributed" *)
logic [WIDTH-1:0] mem [MAX_DEPTH-1:0];
logic [7:0] ptr;

always_ff @(posedge clk) begin
    if(rst) begin
        dout <= '0;
        ptr <= '0;
    end else if(en) begin
        if(delay_depth <= 1) begin
            // Bypass memory: just a register = 1 cycle delay
            dout <= din;
        end else begin
            // Buffer of (delay_depth-1) entries + registered output = delay_depth total
            dout <= mem[ptr];
            mem[ptr] <= din;

            if(ptr >= delay_depth - 2) ptr <= '0;
            else ptr <= ptr + 1'b1;
        end
    end
end

endmodule
